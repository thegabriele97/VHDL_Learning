pll_altera_inst : pll_altera PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
